`timescale 1ns / 10ps

module tx_phy_manager #(
    
) (
    input logic clk, n_rst,

);





endmodule