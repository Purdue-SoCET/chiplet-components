`timescale 1ns / 10ps

module .o #(
    // parameters
) (
    input clk, n_rst
);



endmodule

