`timescale 1ns / 10ps

module tx_phy_manager #() (
    input logic clk, n_rst,
    phy_manager_if.tx_phy phy_if,
    phy_manager_if.tx_switch switch_if
);
    always_comb begin //8b10b encode
        




    end

endmodule