`timescale 1ns / 10ps

module switch #(
    
) (
    input logic clk, n_rst,

);





endmodule