`timescale 1ns / 10ps

module dec_8b10b #(
    // parameters
) (
    input clk, n_rst
);



endmodule

