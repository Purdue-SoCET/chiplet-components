`timescale 1ns / 10ps

module rx_phy_manager #(
    
) (
    input logic clk, n_rst,

);





endmodule