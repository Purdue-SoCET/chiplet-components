
`ifndef SWITCH_VH
`define SWITCH_VH

`include "chiplet_types_pkg.vh"

interface switch_if

    import chiplet_types_pkg::*;

    

    

endinterface

`endif //SWITCH_VH