`include "chiplet_types_pkg.vh"

module cache#(
    parameter NUM_WORDS=128,
    parameter RX = 0
)(
    input logic clk, n_rst,
    input flit_t in_flit,
    input logic data_ready,
    bus_protocol_if.peripheral_vital bus_if
);
    import chiplet_types_pkg::*;

    localparam ADDR_LEN = $clog2(NUM_WORDS);

    logic [31:0] rx_addr, next_rx_addr;
    

    word_t byte_en;

    // TODO: SRAM?
    word_t [NUM_WORDS-1:0] cache, next_cache;

    always_ff @(posedge clk, negedge n_rst) begin
        if (!n_rst) begin
            cache <= '0;
            rx_addr <= '0;
        end else begin
            cache <= next_cache;
            rx_addr <= next_rx_addr
        end
    end

    assign bus_if.rdata = bus_if.ren ? cache[bus_if.addr[2+:ADDR_LEN]] : 32'hBAD1BAD1;
    assign bus_if.request_stall = 0;

    // Expand byte_en to 32 bit signal
    always_comb begin
        for (int i = 0; i < 4; i = i + 1) begin
            byte_en[i*8+:8] = bus_if.strobe[i] ? 8'hFF : 8'h00;
        end
    end

    always_comb begin
        next_cache = cache;
        next_rx_addr = rx_addr;
        if (bus_if.wen || data_ready) begin
            if(RX == 1) begin
                next_cache[rx_addr] = in_flit.payload;
                next_rx_addr += rx_addr + 8;
            end else begin 
                next_cache[bus_if.addr[2+:ADDR_LEN]] = bus_if.wdata & byte_en;
            end
        end
    end
endmodule
