`include "chiplet_types_pkg.vh"

module req_fifo#(
    parameter DEPTH = 16
) (
    input logic clk, n_rst,
    input logic crc_valid,
    input node_id_t req,
    output logic overflow,
    bus_protocol_if.peripheral_vital bus_if
);

    localparam COUNT_ADDR = 32'h3400;
    localparam OVERRUN_ADDR = 32'h3404;
    localparam UNDERRUN_ADDR = 32'h3408;
    localparam REN_ADDR = 32'h340C;

    logic ren, underrun, next_overflow;
    node_id_t next_rdata, rdata, fifo_read, count;

    socetlib_fifo #(.T(logic[4:0]), .DEPTH(DEPTH)) requestor_fifo (
        .CLK(clk),
        .nRST(n_rst),
        .WEN(crc_valid),
        .REN(ren),
        .wdata(req),
        .clear(0),
        .full(),
        .empty(),
        .underrun(underrun),
        .overrun(overflow),
        .count(count),
        .rdata(fifo_read)
    );

always_ff @(posedge clk, negedge n_rst) begin
    if(!n_rst) begin
        rdata <= '0;
    end 
    else begin
        rdata <= next_rdata;
    end
end

always_comb begin
    next_rdata = '0;
    ren = 0;

    if(bus_if.ren) begin
        casez(bus_if.addr)
            COUNT_ADDR: begin
                next_rdata = count;
            end
            OVERRUN_ADDR: begin
                next_rdata = overflow;
            end
            UNDERRUN_ADDR: begin
                next_rdata = underrun;
            end
            REN_ADDR: begin
                ren = 1'b1;
                next_rdata = fifo_read;
            end
            default : begin end
        endcase
    end
end


endmodule
